parameter PATH_WIDTH = <path_width>;
parameter RADIX_WIDTH = <radix_width>;