package lut_pkg;
    localparam TABLE_SIZE = <table_size>;
    localparam SHIFT_VAL = <shift_val>;
    localparam signed MAX_VAL = <max_val>;
    localparam signed MIN_VAL = <min_val>;
endpackage