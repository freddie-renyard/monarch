package tile_pkg;
    localparam SHIFT_VAL = <shift_val>;
    localparam MAX_VAL = <max_val>;
    localparam MIN_VAL = <min_val>;
endpackage