package lut_float_pkg;
    localparam MAN_TABLE_SIZE = <man_table_size>;
    localparam EXP_TABLE_SIZE = <exp_table_size>;
endpackage